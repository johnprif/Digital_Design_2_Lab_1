library verilog;
use verilog.vl_types.all;
entity dec_2_4_vlg_vec_tst is
end dec_2_4_vlg_vec_tst;
