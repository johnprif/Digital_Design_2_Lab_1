library verilog;
use verilog.vl_types.all;
entity my_tff_vlg_vec_tst is
end my_tff_vlg_vec_tst;
