library verilog;
use verilog.vl_types.all;
entity dec_2_4_vlg_check_tst is
    port(
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dec_2_4_vlg_check_tst;
