library verilog;
use verilog.vl_types.all;
entity MyFirstProject_vlg_vec_tst is
end MyFirstProject_vlg_vec_tst;
