library verilog;
use verilog.vl_types.all;
entity my_jkff_vlg_vec_tst is
end my_jkff_vlg_vec_tst;
